package parameter_pkg;
	parameter DATA_WIDTH = 8;
	parameter DEPTH 	 = 8;
	parameter ADDR_WIDTH = $clog2(DATA_WIDTH);
endpackage 